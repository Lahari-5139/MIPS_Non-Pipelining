module instruction_memory(clk,pc, instruction);

input clk;
input[31:0] pc;
output[31:0] instruction;
reg[31:0] instruction;

//256 registers of 32-bits each
reg[31:0] instr_memory[255:0]; 


//MIPS assembly program in binary format
initial 
begin

//LW instructions
instr_memory[0] = 32'b10001100000000010000000000000000;
instr_memory[1] = 32'b10001100000000100000000000000001;
instr_memory[2] = 32'b10001100000000110000000000000010;
instr_memory[3] = 32'b10001100000001000000000000000011;
instr_memory[4] = 32'b10001100000001010000000000000100;
instr_memory[5] = 32'b10001100000001100000000000000101;
instr_memory[6] = 32'b10001100000001110000000000000110;
instr_memory[7] = 32'b10001100000010000000000000000111;
instr_memory[8] = 32'b00000000001001010101000000100001;

//MULT and ADD instructions
instr_memory[9] = 32'b00000000001001010101000000100001; //1 and 5 to 10
instr_memory[10] = 32'b00000000010001110101100000100001; // 2 and 7 to 11
instr_memory[11] = 32'b00000000011001010110000000100001; // 3 and 5 to 12
instr_memory[12] = 32'b00000000100001110110100000100001; // 4 and 7 to 13
instr_memory[13] = 32'b00000000001001100111000000100001; //1 and 6 to 14
instr_memory[14] = 32'b00000000010010000111100000100001; // 2 and 8 to 15
instr_memory[15] = 32'b00000000011001101000000000100001; // 3 and 6 to 16
instr_memory[16] = 32'b00000000100010001000100000100001; // 4 and 8 to 17

//Output Matrix
instr_memory[17] = 32'b00000001010010111010000000100000; // 10 + 11 = 20
instr_memory[18] = 32'b00000001110011111010100000100000; // 14 + 15 = 21
instr_memory[19] = 32'b00000001100011011011000000100000; // 12 + 13 = 33
instr_memory[20] = 32'b00000010000100011011100000100000; // 16 + 17 = 23


end


//Instruction fetch
always @(*)
begin
    instruction = instr_memory[pc];
end

endmodule
