module instruction_memory(clk,pc, instruction);

input clk;
input[31:0] pc;
output[31:0] instruction;
reg[31:0] instruction;

//256 registers of 32-bits each
reg[31:0] instr_memory[255:0]; 


//MIPS assembly program in binary format
initial 
begin

//LW instructions
instr_memory[0] = 32'b10001100000000010000000000000000;
instr_memory[1] = 32'b10001100000000100000000000000001;
instr_memory[2] = 32'b10001100000000110000000000000010;
instr_memory[3] = 32'b10001100000001000000000000000011;
instr_memory[4] = 32'b10001100000001010000000000000100;
instr_memory[5] = 32'b10001100000001100000000000000101;
instr_memory[6] = 32'b10001100000001110000000000000110;
instr_memory[7] = 32'b10001100000010000000000000000111;
instr_memory[8] = 32'b00000000001001010101000000100001;

//MULT and ADD instructions
instr_memory[9] = 32'b00000000001001010101000000100001; //1 and 5 to 10
instr_memory[10] = 32'b00000000010001110101100000100001; // 2 and 7 to 11
instr_memory[11] = 32'b00000000011001010110000000100001; // 3 and 5 to 12
instr_memory[12] = 32'b00000000100001110110100000100001; // 4 and 7 to 13
instr_memory[13] = 32'b00000000001001100111000000100001; //1 and 6 to 14
instr_memory[14] = 32'b00000000010010000111100000100001; // 2 and 8 to 15
instr_memory[15] = 32'b00000000011001101000000000100001; // 3 and 6 to 16
instr_memory[16] = 32'b00000000100010001000100000100001; // 4 and 8 to 17

//Output Matrix
instr_memory[17] = 32'b00000001010010111010000000100000; // 10 + 11 = 20
instr_memory[18] = 32'b00000001110011111010100000100000; // 14 + 15 = 21
instr_memory[19] = 32'b00000001100011011011000000100000; // 12 + 13 = 33
instr_memory[20] = 32'b00000010000100011011100000100000; // 16 + 17 = 23


//instr_memory[0] <= 32'b10001100000000000000000000000000
//instr_memory[1] <= 32'b10001100000000100000000000000010;
//instr_memory[2] <= 32'b10001100000000110000000000110000;
// instr_memory[8] <= 32'b10001100000010010000000000001000;
// instr_memory[9] <= 32'b10001100000010100000000000001001;
// instr_memory[10] <= 32'b10001100000010110000000000001010;
// instr_memory[11] <= 32'b10001100000011000000000000001011;
// instr_memory[12] <= 32'b10001100000011010000000000001100;
// instr_memory[13] <= 32'b10001100000011100000000000001101;
// instr_memory[14] <= 32'b10001100000011110000000000001110;
// instr_memory[15] <= 32'b10001100000100000000000000001111;
// instr_memory[16] <= 32'b10001100000100010000000000010000;
// instr_memory[17] <= 32'b10001100000100100000000000010001;
// instr_memory[12] <= 32'b00000001001010101010000000100000; 
// instr_memory[13] <= 32'b00000000010011011010100000100001;
// instr_memory[20] <= 32'b00000000011100001111000000100001;
// instr_memory[11] <= 32'b00000001001010100101100000100000;
// instr_memory[22] <= 32'b00000011101111101110000000100000;
// instr_memory[23] <= 32'b10101100000100110000000000011100;
// //C01;
// instr_memory[24] <= 32'b00000000001010110000000000100001;
// instr_memory[25] <= 32'b00000000010011101111100000100001;
// instr_memory[26] <= 32'b00000000011100011111000000100001;
// instr_memory[27] <= 32'b00000000000111111110100000100000;
// instr_memory[28] <= 32'b00000011101111101110000000100000;
// instr_memory[29] <= 32'b10101100000101000000000000011100;
// //C02;<
// instr_memory[30] <= 32'b00000000001011000000000000100001;
// instr_memory[31] <= 32'b00000000010011111111100000100001;
// instr_memory[32] <= 32'b00000000011100101111000000100001;
// instr_memory[33] <= 32'b00000000000111111110100000100000;
// instr_memory[34] <= 32'b00000011101111101110000000100000;
// instr_memory[35] <= 32'b10101100000101010000000000011100;
// //C10;<
// instr_memory[36] <= 32'b00000000100010100000000000100001;
// instr_memory[37] <= 32'b00000000101011011111100000100001;
// instr_memory[38] <= 32'b00000000110100001111000000100001;
// instr_memory[39] <= 32'b00000000000111111110100000100000;
// instr_memory[40] <= 32'b00000011101111101110000000100000;
// instr_memory[41] <= 32'b10101100000101100000000000011100;
// //C11;<
// instr_memory[42] <= 32'b00000000100010110000000000100001;
// instr_memory[43] <= 32'b00000000101011101111100000100001;
// instr_memory[44] <= 32'b00000000110100011111000000100001;
// instr_memory[45] <= 32'b00000000000111111110100000100000;
// instr_memory[46] <= 32'b00000011101111101110000000100000;
// instr_memory[47] <= 32'b10101100000101110000000000011100;
// //C12<
// instr_memory[48] <= 32'b00000000100011000000000000100001;
// instr_memory[49] <= 32'b00000000101011111111100000100001;
// instr_memory[50] <= 32'b00000000110100101111000000100001;
// instr_memory[51] <= 32'b00000000000111111110100000100000;
// instr_memory[52] <= 32'b00000011101111101110000000100000;
// instr_memory[53] <= 32'b10101100000110000000000000011100;
// //C20<
// instr_memory[54] <= 32'b00000000111010100000000000100001;
// instr_memory[55] <= 32'b00000001000011011111100000100001;
// instr_memory[56] <= 32'b00000001001100001111000000100001;
// instr_memory[57] <= 32'b00000000000111111110100000100000;
// instr_memory[58] <= 32'b00000011101111101110000000100000;
// instr_memory[59] <= 32'b10101100000110010000000000011100;
// //C21<
// instr_memory[60] <= 32'b00000000111010110000000000100001;
// instr_memory[61] <= 32'b00000001000011101111100000100001;
// instr_memory[62] <= 32'b00000001001100011111000000100001;
// instr_memory[63] <= 32'b00000000000111111110100000100000;
// instr_memory[64] <= 32'b00000011101111101110000000100000;
// instr_memory[65] <= 32'b10101100000110100000000000011100;
// //C22<
// instr_memory[66] <= 32'b00000000111010100000000000100001;
// instr_memory[67] <= 32'b00000001000011111111100000100001;
// instr_memory[68] <= 32'b00000001001100101111000000100001;
// instr_memory[69] <= 32'b00000000000111111110100000100000;
// instr_memory[70] <= 32'b00000011101111101110000000100000;
// instr_memory[71] <= 32'b10101100000110110000000000011100;
end


//Instruction fetch
always @(*)
begin
    instruction = instr_memory[pc];
end

endmodule
